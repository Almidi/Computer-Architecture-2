library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
entity ReorderBuffer is
	Port (
		
		);
end ReorderBuffer;
architecture Structural of ReorderBuffer is
begin
end Structural;